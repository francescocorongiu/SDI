LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Rom_async IS
PORT       (ADDR            : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				OUTPUT         : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END Rom_async;

ARCHITECTURE Behavior OF Rom_async IS
type Rom_type is array (0 to 18) of std_logic_vector(31 downto 0);

constant rom: Rom_type:=(  "00000010000001100000000000000000", --19 elementi della rom da 32 bit ciascuno
									"00000001000001100000000000000000",
									"00000000110001001000000000000000",
									"00000000011000011000000000000000",
									"00000000010000011010000000000000",
									"00000000011000001011000010000000",
									"10110100000000000110001100000000",
									"00000000001010000111110111110000",
									"00000000000000000000000011111000",
									"00000000000000000000100100110110",
									"00000000000000000000000001111001",
									"00000000000000000000000000100110",
									"00000000000000000000000000000000",
									"00000000001011100111110111110000",
									"00000001110001001000000011111000",
									"00000000011000011000100100110110",
									"00000000010000011010000001111001",
									"00000000011000001011000010100110",
									"10110100000000000110001100000000"
									);

BEGIN

 OUTPUT<=rom(to_integer(unsigned(ADDR)));


END Behavior;